`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_2_1 # (parameter N = 4)(

    input [N-1:0] A,
    input [N-1:0] B, 
    input sel,
    output [N-1:0]Y
    );
    
    assign Y = (sel == 1'b1)? B:A;
    
endmodule
